module mux16n1([15:0]a,[3:0]s,[3:0]y,z);
  input[15:0],[3:0]
