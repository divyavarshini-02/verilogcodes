module new(y,a);
output [5:0]y;
input [2:0]a;
assign y=a*a;
endmodule


