module switch_led ()