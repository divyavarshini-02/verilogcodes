`define FPGA_OR_SIMULATION
//`define ASIC_SYNTH
