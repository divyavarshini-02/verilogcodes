/*-------------------------------------------------------------------------------------------------------------------
Design Name : Finite State Machine in a mealy model for 101101 which is overlapping
File name : mealy_1001.v
Desigmer Name: VK. Divyavarshini & S.Santhosh
-------------------------------------------------------------------------------------------------------------------*/
module mealy_101101 ( 
    clk     , //clock
    rst_n   , //syn active low reset
    in      , //input
    out     , //output
);

//----------------------------------------- INPUT PORTS ------------------------------------------------------------//

input clk, rst_n, in;

//----------------------------------------- OUTPUT PORTS -----------------------------------------------------------//

output out;

//----------------------------------------- INPUT DATA TYPES -------------------------------------------------------//

wire in;

//----------------------------------------- OUTPUT DATA TYPES ------------------------------------------------------//

reg out;