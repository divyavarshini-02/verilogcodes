module crc_32(ploy,data,out);
  input [32:0] ploy=33'h104c11db7;
  input [479:0]data;
  output out;

