module top_module()
