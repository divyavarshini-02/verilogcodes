module  ms_7seg_decoder_out()