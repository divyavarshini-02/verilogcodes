module clk(enable,clk_out);
input enable;
output reg clk_out;
