/*-------------------------------------------------------------------------------------------------------------------
Design Name : Finite State Machine in a mealy and moore model for 101 
File name :   MEALY_MOORE_101.v
-------------------------------------------------------------------------------------------------------------------*/
module MEALY_MOORE_101(
);
//----------------------------------------- INPUT PORTS ------------------------------------------------------------//
//----------------------------------------- OUTPUT PORTS -----------------------------------------------------------//
//----------------------------------------- INPUT DATA TYPES -------------------------------------------------------//
//----------------------------------------- OUTPUT DATA TYPES ------------------------------------------------------//
//----------------------------------------- INTERNAL CONSTANTS -----------------------------------------------------//
//----------------------------------------- INTERNAL VARIABLES -----------------------------------------------------//
//----------------------------------------- COMBINATIONAL LOGIC ----------------------------------------------------//
//----------------------------------------- SEQUENTIAL LOGIC -------------------------------------------------------//
//----------------------------------------- OUTPUT LOGIC -----------------------------------------------------------//

endmodule