module name();
reg[795:0]mem[92:0];


integer		var,fd;

initial
begin   
mem[0]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[1]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[2]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[3]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[4]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111100000000001111111111111111111111111111111111111000000011111111111111111111110000000011111111111111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[5]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111110000000000000000000000000000011111111111111111111111111111111111000000000000011111111111111111111111111111111110000000001111111111111111111100000000001111111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111111111110000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[6]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111000000000000000000000000000000000111111111111111111111111111111110000000000000001111111111111111111111111111111110000000001111111111111111111100000000001111111111111111111111111111111111000000000000000000000000000000011111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[7]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111100000000000000000000000000000000000001111111111111111111111111111110000000000000000111111111111111111111111111111110000000001111111111111111111100000000001111111111111111111111111111111100000000000000000000000000000000001111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[8]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111110000000000000000000000000000000000000000011111111111111111111111111110000000000000000011111111111111111111111111111110000000001111111111111111111100000000001111111111111111111111111111111000000000000000000000000000000000000011111111111111111111111111111111100000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[9]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111100000000000000000000000000000000000000000001111111111111111111111111110000000000000000011111111111111111111111111111110000000001111111111111111111100000000001111111111111111111111111111100000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[10]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011111111111111111111111111111111111111111111100000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111110000000000000000001111111111111111111111111111110000000001111111111111111111100000000001111111111111111111111111111000000000000000000000000000000000000000000111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[11]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111100000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000011111111111111111111111110000000000000000001111111111111111111111111111110000000001111111111111111111100000000001111111111111111111111111110000000000000000000000000000000000000000000111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[12]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111000000000000000000001111111111111111111111111100000000000000001111111111111111000000000000000001111111111111111111111110000000000000000000111111111111111111111111111110000000001111111111111111111100000000001111111111111111111111111100000000000000000111111111111100000000000000111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[13]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111000000000100000000001111111111111111111111111000000000000000111111111111111111110000000000000000111111111111111111111110000000000000000000111111111111111111111111111110000000001111111111111111111100000000001111111111111111111111111000000000000000111111111111111111100000000000111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[14]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000010000000000111111111111111111111111111111111111111111000000000100000000001111111111111111111111110000000000000011111111111111111111111100000000000000011111111111111111111110000000000000000000011111111111111111111111111110000000001111111111111111111100000000001111111111111111111111110000000000000011111111111111111111111000000000111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[15]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000010000000000111111111111111111111111111111111111111110000000001100000000001111111111111111111111100000000000000111111111111111111111111111000000000000011111111111111111111110000000000000000000001111111111111111111111111110000000001111111111111111111100000000001111111111111111111111100000000000000111111111111111111111111110000000111111111111111111111111111110000000001000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[16]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011000000000011111111111111111111111111111111111111110000000001100000000001111111111111111111111000000000000011111111111111111111111111111100000000000001111111111111111111110000000000000000000001111111111111111111111111110000000001111111111111111111100000000001111111111111111111111100000000000001111111111111111111111111111100000111111111111111111111111111100000000011000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[17]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011000000000011111111111111111111111111111111111111100000000001100000000001111111111111111111111000000000000111111111111111111111111111111110000000000000111111111111111111110000000000100000000000111111111111111111111111110000000001111111111111111111100000000001111111111111111111111000000000000011111111111111111111111111111110000111111111111111111111111111100000000011100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[18]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011000000000011111111111111111111111111111111111111100000000011100000000001111111111111111111110000000000001111111111111111111111111111111111000000000000111111111111111111110000000000100000000000111111111111111111111111110000000001111111111111111111100000000001111111111111111111111000000000000111111111111111111111111111111111101111111111111111111111111111100000000011100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[19]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011100000000001111111111111111111111111111111111111000000000011100000000001111111111111111111110000000000001111111111111111111111111111111111100000000000011111111111111111110000000000110000000000011111111111111111111111110000000001111111111111111111100000000001111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111000000000111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[20]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011100000000001111111111111111111111111111111111111000000000111100000000001111111111111111111100000000000011111111111111111111111111111111111100000000000011111111111111111110000000000110000000000011111111111111111111111110000000001111111111111111111100000000001111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111000000000111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[21]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011110000000000111111111111111111111111111111111111000000000111100000000001111111111111111111100000000000111111111111111111111111111111111111110000000000001111111111111111110000000000111000000000001111111111111111111111110000000001111111111111111111100000000001111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111110000000000111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[22]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011110000000000111111111111111111111111111111111110000000000111100000000001111111111111111111000000000000111111111111111111111111111111111111110000000000001111111111111111110000000000111000000000001111111111111111111111110000000001111111111111111111100000000001111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111110000000001111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[24]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011110000000000011111111111111111111111111111111110000000001111100000000001111111111111111111000000000001111111111111111111111111111111111111111000000000001111111111111111110000000000111100000000000111111111111111111111110000000001111111111111111111100000000001111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111110000000001111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[25]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111000000000011111111111111111111111111111111100000000001111100000000001111111111111111111000000000001111111111111111111111111111111111111111000000000000111111111111111110000000000111100000000000011111111111111111111110000000001111111111111111111100000000001111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111100000000001111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[26]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111000000000011111111111111111111111111111111100000000011111100000000001111111111111111110000000000011111111111111111111111111111111111111111100000000000111111111111111110000000000111110000000000011111111111111111111110000000001111111111111111111100000000001111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111100000000011111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[27]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111100000000001111111111111111111111111111111000000000011111100000000001111111111111111110000000000011111111111111111111111111111111111111111100000000000111111111111111110000000000111110000000000001111111111111111111110000000001111111111111111111100000000001111111111111111110000000000011111111111111111111111111111111111111111111111111111111111111111100000000011111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[28]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111100000000001111111111111111111111111111111000000000111111100000000001111111111111111110000000000111111111111111111111111111111111111111111100000000000111111111111111110000000000111111000000000001111111111111111111110000000001111111111111111111100000000001111111111111111110000000000011111111111111111111111111111111111111111111111111111111111111111000000000011111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[29]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111100000000000111111111111111111111111111111000000000111111100000000001111111111111111100000000000111111111111111111111111111111111111111111110000000000011111111111111110000000000111111000000000000111111111111111111110000000001111111111111111111100000000001111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111000000000111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[30]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111110000000000111111111111111111111111111110000000000111111100000000001111111111111111100000000000111111111111111111111111111111111111111111110000000000011111111111111110000000000111111100000000000111111111111111111110000000001111111111111111111100000000001111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111000000000111111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[31]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111110000000000111111111111111111111111111110000000001111111100000000001111111111111111100000000000111111111111111111111111111111111111111111110000000000011111111111111110000000000111111110000000000011111111111111111110000000001111111111111111111100000000001111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111110000000000111111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[32]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111000000000011111111111111111111111111100000000001111111100000000001111111111111111100000000001111111111111111111111111111111111111111111110000000000011111111111111110000000000111111110000000000011111111111111111110000000001111111111111111111100000000001111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111110000000001111111111110000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[33]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111000000000011111111111111111111111111100000000011111111100000000001111111111111111100000000001111111111111111111111111111111111111111111110000000000011111111111111110000000000111111111000000000001111111111111111110000000001111111111111111111100000000001111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111100000000001111111111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[34]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111000000000001111111111111111111111111100000000011111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000011111111111111110000000000111111111000000000000111111111111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111100000000001111111111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[35]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111100000000001111111111111111111111111000000000011111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000011111111111111110000000000111111111100000000000111111111111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111100000000011111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[36]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111100000000001111111111111111111111111000000000111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000011111111111111110000000000111111111100000000000011111111111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111000000000011111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[37]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111100000000000111111111111111111111110000000000111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000001111111111111110000000000111111111110000000000011111111111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111000000000011111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[38]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111110000000000111111111111111111111110000000001111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000001111111111111110000000000111111111111000000000001111111111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111000000000111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[39]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111110000000000011111111111111111111100000000001111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000001111111111111110000000000111111111111000000000001111111111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111111110000000000111111111111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[40]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111000000000011111111111111111111100000000001111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000001111111111111110000000000111111111111100000000000111111111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111111110000000001111111111111111110000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[41]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111000000000011111111111111111111100000000011111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000001111111111111110000000000111111111111100000000000111111111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111111110000000001111111111111111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[42]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111000000000001111111111111111111000000000011111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000001111111111111110000000000111111111111110000000000011111111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111111100000000001111111111111111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[43]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111100000000001111111111111111111000000000111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000001111111111111110000000000111111111111110000000000011111111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[44]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111100000000000111111111111111110000000000111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000001111111111111110000000000111111111111111000000000001111111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[45]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111110000000000111111111111111110000000000111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000001111111111111110000000000111111111111111000000000000111111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[46]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111110000000000111111111111111110000000001111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000001111111111111110000000000111111111111111100000000000111111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[47]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111110000000000011111111111111100000000001111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000011111111111111110000000000111111111111111110000000000011111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[48]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111000000000011111111111111100000000011111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000011111111111111110000000000111111111111111110000000000011111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111110000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[49]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111000000000001111111111111000000000011111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000011111111111111110000000000111111111111111111000000000001111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111110000000001111111111111111111111110000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[50]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111100000000001111111111111000000000011111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111000000000011111111111111110000000000111111111111111111000000000001111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111100000000001111111111111111111111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[51]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111100000000001111111111110000000000111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111110000000000011111111111111110000000000111111111111111111100000000000111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111100000000001111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[52]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111100000000000111111111110000000000111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111110000000000011111111111111110000000000111111111111111111100000000000111111110000000001111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[53]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111110000000000111111111110000000001111111111111111100000000001111111111111111100000000001111111111111111111111111111111111111111111110000000000011111111111111110000000000111111111111111111110000000000011111110000000001111111111111111111100000000001111111111111111000000000000111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[54]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111110000000000011111111100000000001111111111111111100000000001111111111111111100000000000111111111111111111111111111111111111111111110000000000011111111111111110000000000111111111111111111110000000000001111110000000001111111111111111111100000000001111111111111111100000000000111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[55]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111000000000011111111100000000011111111111111111100000000001111111111111111100000000000111111111111111111111111111111111111111111110000000000111111111111111110000000000111111111111111111111000000000001111110000000001111111111111111111100000000001111111111111111100000000000111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[56]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111000000000011111111000000000011111111111111111100000000001111111111111111100000000000111111111111111111111111111111111111111111100000000000111111111111111110000000000111111111111111111111100000000000111110000000001111111111111111111100000000001111111111111111100000000000111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[57]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111000000000001111111000000000011111111111111111100000000001111111111111111100000000000111111111111111111111111111111111111111111100000000000111111111111111110000000000111111111111111111111100000000000111110000000001111111111111111111100000000001111111111111111100000000000011111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[58]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111100000000001111111000000000111111111111111111100000000001111111111111111100000000000011111111111111111111111111111111111111111100000000000111111111111111110000000000111111111111111111111110000000000011110000000001111111111111111111100000000001111111111111111100000000000011111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[59]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111100000000000111110000000000111111111111111111100000000001111111111111111110000000000011111111111111111111111111111111111111111000000000001111111111111111110000000000111111111111111111111110000000000011110000000001111111111111111111100000000001111111111111111110000000000011111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[60]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111100000000000111110000000001111111111111111111100000000001111111111111111110000000000011111111111111111111111111111111111111111000000000001111111111111111110000000000111111111111111111111111000000000001110000000001111111111111111111100000000001111111111111111110000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[61]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111110000000000111100000000001111111111111111111100000000001111111111111111110000000000001111111111111111111111111111111111111110000000000001111111111111111110000000000111111111111111111111111000000000001110000000001111111111111111111100000000001111111111111111110000000000001111111111111111111111111111111111111111111111111111000000000011111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[62]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111110000000000011100000000001111111111111111111100000000001111111111111111111000000000001111111111111111111111111111111111111110000000000011111111111111111110000000000111111111111111111111111100000000000110000000001111111111111111111100000000001111111111111111111000000000000111111111111111111111111111111111111111111111111111000000000011111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[63]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111000000000011000000000011111111111111111111100000000001111111111111111111000000000000111111111111111111111111111111111111100000000000011111111111111111110000000000111111111111111111111111100000000000110000000001111111111111111111100000000001111111111111111111000000000000111111111111111111111111111111111111111111111111111000000000011111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[64]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111000000000001000000000011111111111111111111100000000001111111111111111111000000000000111111111111111111111111111111111111100000000000111111111111111111110000000000111111111111111111111111110000000000010000000001111111111111111111100000000001111111111111111111100000000000011111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[65]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111000000000001000000000111111111111111111111100000000001111111111111111111100000000000011111111111111111111111111111111111000000000000111111111111111111110000000000111111111111111111111111111000000000010000000001111111111111111111100000000001111111111111111111100000000000001111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[66]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111100000000000000000000111111111111111111111100000000001111111111111111111100000000000001111111111111111111111111111111110000000000001111111111111111111110000000000111111111111111111111111111000000000000000000001111111111111111111100000000001111111111111111111110000000000000111111111111111111111111111111111100111111111100000000000111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[67]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111100000000000000000000111111111111111111111100000000001111111111111111111110000000000000111111111111111111111111111111100000000000001111111111111111111110000000000111111111111111111111111111100000000000000000001111111111111111111100000000001111111111111111111110000000000000011111111111111111111111111111110000011111111100000000001111111111111111111111111111111111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[68]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111110000000000000000001111111111111111111111100000000001111111111111111111110000000000000011111111111111111111111111111000000000000011111111111111111111110000000000111111111111111111111111111100000000000000000001111111111111111111100000000001111111111111111111111000000000000001111111111111111111111111111100000011111111100000000001111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[69]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111110000000000000000001111111111111111111111100000000001111111111111111111111000000000000001111111111111111111111111110000000000000111111111111111111111110000000000111111111111111111111111111110000000000000000001111111111111111111100000000001111111111111111111111000000000000000111111111111111111111111110000000011111111000000000001111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[70]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111110000000000000000011111111111111111111111100000000001111111111111111111111100000000000000111111111111111111111111000000000000000111111111111111111111110000000000111111111111111111111111111110000000000000000001111111111111111111100000000001111111111111111111111100000000000000011111111111111111111111000000000011111111000000000011111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[71]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111000000000000000011111111111111111111111100000000001111111111111111111111100000000000000000111111111111111111100000000000000001111111111111111111111110000000000111111111111111111111111111111000000000000000001111111111111111111100000000001111111111111111111111110000000000000000011111111111111111100000000000011111111000000000011111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[72]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111000000000000000011111111111111111111111100000000001111111111111111111111110000000000000000001111111111111100000000000000000011111111111111111111111110000000000111111111111111111111111111111000000000000000001111111111111111111100000000001111111111111111111111111000000000000000000011111111111000000000000000011111110000000000011111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[73]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111100000000000000111111111111111111111111100000000001111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111110000000000111111111111111111111111111111100000000000000001111111111111111111100000000001111111111111111111111111100000000000000000000000000000000000000000000111111110000000000111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[74]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111100000000000000111111111111111111111111100000000001111111111111111111111111100000000000000000000000000000000000000000000001111111111111111111111111110000000000111111111111111111111111111111110000000000000001111111111111111111100000000001111111111111111111111111110000000000000000000000000000000000000000000111111110000000000111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[75]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111100000000000001111111111111111111111111100000000001111111111111111111111111110000000000000000000000000000000000000000000011111111111111111111111111110000000000111111111111111111111111111111110000000000000001111111111111111111100000000001111111111111111111111111111000000000000000000000000000000000000000001111111100000000000111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[76]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111110000000000001111111111111111111111111100000000001111111111111111111111111111100000000000000000000000000000000000000001111111111111111111111111111110000000000111111111111111111111111111111111000000000000001111111111111111111100000000001111111111111111111111111111100000000000000000000000000000000000000111111111100000000001111111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[77]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111110000000000011111111111111111111111111100000000001111111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111111110000000000111111111111111111111111111111111000000000000001111111111111111111100000000001111111111111111111111111111111000000000000000000000000000000000001111111111100000000001111111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[78]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111110000000000011111111111111111111111111100000000001111111111111111111111111111111100000000000000000000000000000000001111111111111111111111111111111110000000000111111111111111111111111111111111100000000000001111111111111111111100000000001111111111111111111111111111111100000000000000000000000000000000111111111111000000000001111111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[79]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111111000000000011111111111111111111111111100000000001111111111111111111111111111111111000000000000000000000000000001111111111111111111111111111111111110000000000111111111111111111111111111111111110000000000001111111111111111111100000000001111111111111111111111111111111111100000000000000000000000000111111111111111000000000011111111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[80]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000111111111111111111111111111100000001111111111111111111111111111110000000111111111111111111111111111111111111111000000000000000000000001111111111111111111111111111111111111111000000011111111111111111111111111111111111111100000000111111111111111111111110000000011111111111111111111111111111111111111000000000000000000000111111111111111111100000000111111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[81]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[82]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[83]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[84]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[85]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[86]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[87]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[88]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[89]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[90]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[91]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[92]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[93]=795'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
end



initial
begin
   // $writememb("name_display.bin",mem);
	fd=$fopen("name_display.bin","w");	

	for(var=0;var<93;var=var+1)
	begin
		$fdisplayb(fd,mem[var]);
	end

end
endmodule





