module divyavarshini();
reg[325:0]mem[84:1];
integer fd;

initial
begin

mem[0] = 326'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[1] = 326'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[2] = 326'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[3] = 326'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[4] = 326'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[5] = 326'b1111111111111111111111111111100000000000000000000000000011111111111111111111111111111111111111111111110000000011111111111111000000000111111111111111111111111111111111111111111111000000001111110000000011111111111111111111111111111111111100000000011111111111111111111111111111111000000000011111111111111111111111111111111;
mem[6] = 326'b1111111111111111111111111111000000000000000000000000000000000111111111111111111111111111111111111111100000000001111111111110000000000011111111111111111111111111111111111111111110000000000111100000000000111111111111111111111111111111111000000000001111111111111111111111111111100000000000001111111111111111111111111111111;
mem[7] = 326'b1111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111111111111100000000001111111111110000000000011111111111111111111111111111111111111111110000000000111100000000000111111111111111111111111111111111000000000011111111111111111111111111111100000000000000111111111111111111111111111111;
mem[8] = 326'b1111111111111111111111111110000000000000000000000000000000000000000111111111111111111111111111111111100000000001111111111110000000000011111111111111111111111111111111111111111100000000000111110000000000011111111111111111111111111111110000000000011111111111111111111111111111100000000000000111111111111111111111111111111;
mem[9] = 326'b1111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111111100000000001111111111111000000000001111111111111111111111111111111111111111100000000001111110000000000011111111111111111111111111111110000000000011111111111111111111111111111000000000000000111111111111111111111111111111;
mem[10] =326'b1111111111111111111111111110000000000000000000000000000000000000000000011111111111111111111111111111100000000001111111111111000000000001111111111111111111111111111111111111111100000000001111111000000000001111111111111111111111111111100000000000111111111111111111111111111111000000000000000011111111111111111111111111111;
mem[11] =326'b1111111111111111111111111110000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111111100000000001111111111111111111111111111111111111111000000000001111111000000000001111111111111111111111111111100000000001111111111111111111111111111110000000000000000011111111111111111111111111111;
mem[12] =326'b1111111111111111111111111110000000000000000000000000000000000000000000000111111111111111111111111111100000000001111111111111100000000000111111111111111111111111111111111111111000000000011111111100000000000111111111111111111111111111000000000001111111111111111111111111111110000000000000000011111111111111111111111111111;
mem[13] =326'b1111111111111111111111111110000000000111111111111110000000000000000000000001111111111111111111111111100000000001111111111111100000000000111111111111111111111111111111111111111000000000011111111100000000000111111111111111111111111111000000000011111111111111111111111111111110000000000000000001111111111111111111111111111;
mem[14] =326'b1111111111111111111111111110000000000111111111111111111110000000000000000000111111111111111111111111100000000001111111111111110000000000111111111111111111111111111111111111110000000000011111111110000000000011111111111111111111111110000000000011111111111111111111111111111100000000000000000001111111111111111111111111111;
mem[15] =326'b1111111111111111111111111110000000000111111111111111111111110000000000000000011111111111111111111111100000000001111111111111110000000000011111111111111111111111111111111111110000000000111111111110000000000011111111111111111111111110000000000111111111111111111111111111111100000000000000000000111111111111111111111111111;
mem[16] =326'b1111111111111111111111111110000000000111111111111111111111111111000000000000001111111111111111111111100000000001111111111111111000000000011111111111111111111111111111111111100000000000111111111111000000000001111111111111111111111100000000001111111111111111111111111111111000000000110000000000111111111111111111111111111;
mem[17] =326'b1111111111111111111111111110000000000111111111111111111111111111100000000000000111111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111100000000001111111111111100000000000111111111111111111111000000000001111111111111111111111111111111000000000111000000000011111111111111111111111111;
mem[18] =326'b1111111111111111111111111110000000000111111111111111111111111111110000000000000011111111111111111111100000000001111111111111111000000000001111111111111111111111111111111111100000000001111111111111100000000000111111111111111111111000000000011111111111111111111111111111111000000000111000000000011111111111111111111111111;
mem[19] =326'b1111111111111111111111111110000000000111111111111111111111111111111100000000000011111111111111111111100000000001111111111111111100000000000111111111111111111111111111111111000000000011111111111111110000000000011111111111111111110000000000011111111111111111111111111111110000000001111000000000011111111111111111111111111;
mem[20] =326'b1111111111111111111111111110000000000111111111111111111111111111111100000000000001111111111111111111100000000001111111111111111100000000000111111111111111111111111111111111000000000011111111111111110000000000011111111111111111110000000000111111111111111111111111111111110000000001111100000000001111111111111111111111111;
mem[21] =326'b1111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111100000000001111111111111111100000000000111111111111111111111111111111111000000000011111111111111111000000000001111111111111111100000000000111111111111111111111111111111100000000001111100000000001111111111111111111111111;
mem[22] =326'b1111111111111111111111111110000000000111111111111111111111111111111111000000000000111111111111111111100000000001111111111111111110000000000011111111111111111111111111111110000000000111111111111111111000000000001111111111111111100000000001111111111111111111111111111111100000000011111100000000001111111111111111111111111;
mem[23] =326'b1111111111111111111111111110000000000111111111111111111111111111111111100000000000111111111111111111100000000001111111111111111110000000000011111111111111111111111111111110000000000111111111111111111100000000000111111111111111000000000001111111111111111111111111111111100000000011111110000000000111111111111111111111111;
mem[24] =326'b1111111111111111111111111110000000000111111111111111111111111111111111100000000000011111111111111111100000000001111111111111111110000000000011111111111111111111111111111110000000000111111111111111111100000000000111111111111111000000000011111111111111111111111111111111000000000011111110000000000111111111111111111111111;
mem[25] =326'b1111111111111111111111111110000000000111111111111111111111111111111111110000000000011111111111111111100000000001111111111111111111000000000001111111111111111111111111111100000000001111111111111111111110000000000011111111111110000000000011111111111111111111111111111111000000000111111110000000000011111111111111111111111;
mem[26] =326'b1111111111111111111111111110000000000111111111111111111111111111111111110000000000011111111111111111100000000001111111111111111111000000000001111111111111111111111111111100000000001111111111111111111110000000000011111111111110000000000111111111111111111111111111111111000000000111111111000000000011111111111111111111111;
mem[27] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111000000000001111111111111111100000000001111111111111111111100000000001111111111111111111111111111100000000001111111111111111111111000000000001111111111100000000000111111111111111111111111111111110000000000111111111000000000011111111111111111111111;
mem[28] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111000000000001111111111111111100000000001111111111111111111100000000000111111111111111111111111111000000000011111111111111111111111000000000001111111111100000000001111111111111111111111111111111110000000001111111111000000000001111111111111111111111;
mem[29] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111000000000001111111111111111100000000001111111111111111111100000000000111111111111111111111111111000000000011111111111111111111111100000000001111111111100000000001111111111111111111111111111111110000000001111111111100000000001111111111111111111111;
mem[30] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111100000000001111111111111111100000000001111111111111111111110000000000111111111111111111111111111000000000011111111111111111111111100000000000111111111000000000011111111111111111111111111111111100000000001111111111100000000001111111111111111111111;
mem[31] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111100000000000111111111111111100000000001111111111111111111110000000000011111111111111111111111110000000000111111111111111111111111110000000000111111111000000000011111111111111111111111111111111100000000011111111111100000000000111111111111111111111;
mem[32] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111100000000000111111111111111100000000001111111111111111111110000000000011111111111111111111111110000000000111111111111111111111111110000000000011111110000000000111111111111111111111111111111111000000000011111111111110000000000111111111111111111111;
mem[33] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111100000000000111111111111111100000000001111111111111111111111000000000011111111111111111111111110000000000111111111111111111111111111000000000011111110000000000111111111111111111111111111111111000000000011111111111110000000000111111111111111111111;
mem[34] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111100000000000111111111111111100000000001111111111111111111111000000000001111111111111111111111100000000001111111111111111111111111111000000000001111100000000001111111111111111111111111111111111000000000111111111111110000000000011111111111111111111;
mem[35] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111100000000000111111111111111100000000001111111111111111111111000000000001111111111111111111111100000000001111111111111111111111111111100000000001111100000000001111111111111111111111111111111110000000000111111111111111000000000011111111111111111111;
mem[36] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111110000000000111111111111111100000000001111111111111111111111100000000001111111111111111111111100000000011111111111111111111111111111100000000000111000000000011111111111111111111111111111111110000000000111111111111111000000000001111111111111111111;
mem[37] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111110000000000111111111111111100000000001111111111111111111111100000000000111111111111111111111000000000011111111111111111111111111111110000000000111000000000011111111111111111111111111111111110000000001111111111111111000000000001111111111111111111;
mem[38] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111110000000000111111111111111100000000001111111111111111111111100000000000111111111111111111111000000000011111111111111111111111111111110000000000111000000000111111111111111111111111111111111100000000001111111111111111100000000001111111111111111111;
mem[39] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111110000000000111111111111111100000000001111111111111111111111110000000000111111111111111111111000000000111111111111111111111111111111111000000000010000000000111111111111111111111111111111111100000000011111111111111111100000000000111111111111111111;
mem[40] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111110000000000111111111111111100000000001111111111111111111111110000000000011111111111111111110000000000111111111111111111111111111111111000000000010000000001111111111111111111111111111111111100000000011111111111111111110000000000111111111111111111;
mem[41] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111110000000000111111111111111100000000001111111111111111111111111000000000011111111111111111110000000000111111111111111111111111111111111100000000000000000001111111111111111111111111111111111000000000011111111111111111110000000000111111111111111111;
mem[42] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111110000000000111111111111111100000000001111111111111111111111111000000000011111111111111111110000000001111111111111111111111111111111111100000000000000000011111111111111111111111111111111111000000000111111111111111111110000000000011111111111111111;
mem[43] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111110000000000111111111111111100000000001111111111111111111111111000000000001111111111111111100000000001111111111111111111111111111111111110000000000000000011111111111111111111111111111111110000000000111111111111111111111000000000011111111111111111;
mem[44] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111110000000000111111111111111100000000001111111111111111111111111100000000001111111111111111100000000001111111111111111111111111111111111110000000000000000111111111111111111111111111111111110000000000111111111111111111111000000000011111111111111111;
mem[45] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111110000000000111111111111111100000000001111111111111111111111111100000000001111111111111111100000000011111111111111111111111111111111111111000000000000000111111111111111111111111111111111110000000001111111111111111111111000000000001111111111111111;
mem[46] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111110000000000111111111111111100000000001111111111111111111111111100000000000111111111111111000000000011111111111111111111111111111111111111000000000000001111111111111111111111111111111111100000000001111111111111111111111100000000001111111111111111;
mem[47] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111110000000000111111111111111100000000001111111111111111111111111110000000000111111111111111000000000011111111111111111111111111111111111111100000000000001111111111111111111111111111111111100000000001111111111111111111111100000000000111111111111111;
mem[48] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111100000000000111111111111111100000000001111111111111111111111111110000000000111111111111111000000000111111111111111111111111111111111111111100000000000011111111111111111111111111111111111100000000011111111111111111111111100000000000111111111111111;
mem[49] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111100000000000111111111111111100000000001111111111111111111111111110000000000011111111111110000000000111111111111111111111111111111111111111110000000000011111111111111111111111111111111111000000000011111111111111111111111110000000000111111111111111;
mem[50] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111100000000000111111111111111100000000001111111111111111111111111111000000000011111111111110000000001111111111111111111111111111111111111111110000000000111111111111111111111111111111111111000000000011111111111111111111111110000000000011111111111111;
mem[51] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111100000000000111111111111111100000000001111111111111111111111111111000000000011111111111110000000001111111111111111111111111111111111111111110000000000111111111111111111111111111111111111000000000111111111111111111111111110000000000011111111111111;
mem[52] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111100000000001111111111111111100000000001111111111111111111111111111000000000001111111111100000000001111111111111111111111111111111111111111110000000000111111111111111111111111111111111110000000000000000000000000000000000000000000000011111111111111;
mem[53] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111100000000001111111111111111100000000001111111111111111111111111111100000000001111111111100000000011111111111111111111111111111111111111111110000000000111111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111;
mem[54] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111000000000001111111111111111100000000001111111111111111111111111111100000000000111111111100000000011111111111111111111111111111111111111111110000000000111111111111111111111111111111111100000000000000000000000000000000000000000000000001111111111111;
mem[55] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111000000000001111111111111111100000000001111111111111111111111111111100000000000111111111000000000011111111111111111111111111111111111111111110000000000111111111111111111111111111111111100000000000000000000000000000000000000000000000001111111111111;
mem[56] =326'b1111111111111111111111111110000000000111111111111111111111111111111111111000000000011111111111111111100000000001111111111111111111111111111110000000000111111111000000000111111111111111111111111111111111111111111110000000000111111111111111111111111111111111100000000000000000000000000000000000000000000000000111111111111;
mem[57] =326'b1111111111111111111111111110000000000111111111111111111111111111111111110000000000011111111111111111100000000001111111111111111111111111111110000000000011111111000000000111111111111111111111111111111111111111111110000000000111111111111111111111111111111111000000000000000000000000000000000000000000000000000111111111111;
mem[58] =326'b1111111111111111111111111110000000000111111111111111111111111111111111110000000000011111111111111111100000000001111111111111111111111111111111000000000011111110000000000111111111111111111111111111111111111111111110000000000111111111111111111111111111111111000000000000000000000000000000000000000000000000000011111111111;
mem[59] =326'b1111111111111111111111111110000000000111111111111111111111111111111111100000000000111111111111111111100000000001111111111111111111111111111111000000000011111110000000001111111111111111111111111111111111111111111110000000000111111111111111111111111111111111000000000000000000000000000000000000000000000000000011111111111;
mem[60] =326'b1111111111111111111111111110000000000111111111111111111111111111111111100000000000111111111111111111100000000001111111111111111111111111111111000000000001111110000000001111111111111111111111111111111111111111111110000000000111111111111111111111111111111110000000000111111111111111111111111111111110000000000011111111111;
mem[61] =326'b1111111111111111111111111110000000000111111111111111111111111111111111000000000000111111111111111111100000000001111111111111111111111111111111100000000001111100000000001111111111111111111111111111111111111111111110000000000111111111111111111111111111111110000000000111111111111111111111111111111111000000000001111111111;
mem[62] =326'b1111111111111111111111111110000000000111111111111111111111111111111111000000000001111111111111111111100000000001111111111111111111111111111111100000000001111100000000011111111111111111111111111111111111111111111110000000000111111111111111111111111111111110000000000111111111111111111111111111111111000000000001111111111;
mem[63] =326'b1111111111111111111111111110000000000111111111111111111111111111111110000000000001111111111111111111100000000001111111111111111111111111111111100000000000111100000000011111111111111111111111111111111111111111111110000000000111111111111111111111111111111100000000001111111111111111111111111111111111000000000001111111111;
mem[64] =326'b1111111111111111111111111110000000000111111111111111111111111111111100000000000011111111111111111111100000000001111111111111111111111111111111110000000000111000000000011111111111111111111111111111111111111111111110000000000111111111111111111111111111111100000000001111111111111111111111111111111111100000000000111111111;
mem[65] =326'b1111111111111111111111111110000000000111111111111111111111111111111000000000000111111111111111111111100000000001111111111111111111111111111111110000000000111000000000111111111111111111111111111111111111111111111110000000000111111111111111111111111111111000000000001111111111111111111111111111111111100000000000111111111;
mem[66] =326'b1111111111111111111111111110000000000111111111111111111111111111110000000000000111111111111111111111100000000001111111111111111111111111111111110000000000011000000000111111111111111111111111111111111111111111111110000000000111111111111111111111111111111000000000011111111111111111111111111111111111110000000000111111111;
mem[67] =326'b1111111111111111111111111110000000000111111111111111111111111111000000000000001111111111111111111111100000000001111111111111111111111111111111111000000000010000000001111111111111111111111111111111111111111111111110000000000111111111111111111111111111111000000000011111111111111111111111111111111111110000000000011111111;
mem[68] =326'b1111111111111111111111111110000000000111111111111111111111111110000000000000011111111111111111111111100000000001111111111111111111111111111111111000000000010000000001111111111111111111111111111111111111111111111110000000000111111111111111111111111111110000000000011111111111111111111111111111111111110000000000011111111;
mem[69] =326'b1111111111111111111111111110000000000111111111111111111111111000000000000000111111111111111111111111100000000001111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111110000000000111111111111111111111111111110000000000111111111111111111111111111111111111111000000000001111111;
mem[70] =326'b1111111111111111111111111110000000000111111111111111111111000000000000000001111111111111111111111111100000000001111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111111111110000000000111111111111111111111111111110000000000111111111111111111111111111111111111111000000000001111111;
mem[71] =326'b1111111111111111111111111110000000000111111111111110000000000000000000000011111111111111111111111111100000000001111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111111111110000000000111111111111111111111111111100000000000111111111111111111111111111111111111111000000000001111111;
mem[72] =326'b1111111111111111111111111110000000000000000000000000000000000000000000000111111111111111111111111111100000000001111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111111111110000000000111111111111111111111111111100000000001111111111111111111111111111111111111111100000000000111111;
mem[73] =326'b1111111111111111111111111110000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111110000000000111111111111111111111111111100000000001111111111111111111111111111111111111111100000000000111111;
mem[74] =326'b1111111111111111111111111110000000000000000000000000000000000000000000111111111111111111111111111111100000000001111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111110000000000111111111111111111111111111000000000001111111111111111111111111111111111111111100000000000111111;
mem[75] =326'b1111111111111111111111111110000000000000000000000000000000000000000011111111111111111111111111111111100000000001111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111110000000000111111111111111111111111111000000000011111111111111111111111111111111111111111110000000000011111;
mem[76] =326'b1111111111111111111111111110000000000000000000000000000000000000001111111111111111111111111111111111100000000001111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111110000000000111111111111111111111111111000000000011111111111111111111111111111111111111111110000000000011111;
mem[77] =326'b1111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111111111111100000000001111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111110000000000111111111111111111111111110000000000011111111111111111111111111111111111111111110000000000011111;
mem[78] =326'b1111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111100000000001111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111111111111110000000000111111111111111111111111110000000000111111111111111111111111111111111111111111111000000000011111;
mem[79] =326'b1111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111110000000011111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111111111111000000001111111111111111111111111111000000001111111111111111111111111111111111111111111111100000000011111;
mem[80] =326'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[81] =326'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[82] =326'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[83] =326'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
mem[84] =326'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

end

initial
begin
	fd = $fopen("divyavarshini.bin" ,"w");
end

initial
begin
    $writememb("divyavarshini.bin",mem);
end
endmodule









